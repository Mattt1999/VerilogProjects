module diff(
	input [2:0]a, b,
	output [2:0]out
);

assign out = a - b;

endmodule 