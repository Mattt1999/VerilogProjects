module bitwise_xor(

	input [2:0]a, c,
	output [2:0]out
);

assign out = a ^ c;

endmodule 