module adunare(
	input [1:0]in0, in1,
	output [2:0] out
);

assign out = in0 + in1;

endmodule 