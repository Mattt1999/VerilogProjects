module bitwise_or(
	input [2:0]b, c,
	output [2:0]out

);


assign out = b | c;

endmodule 