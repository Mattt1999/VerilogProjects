module bitwise_not(

	input [2:0]c,
	output [2:0]out

);

assign out = ~c; 

endmodule 